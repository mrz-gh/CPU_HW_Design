module FetchStage (
    clk,
    rst,
    freeze,
    Branch_taken,
    BranchAddr,
    PC,
    Instruction
);
    // parameter INST_NUM = 129;

    input wire clk;
    input wire rst;
    input wire freeze;
    input wire Branch_taken;
    input [31:0] BranchAddr;
    output [31:0] PC;
    output reg [31:0] Instruction;
    
    reg [31:0] PC_Reg;
    wire [31:0] PC_In;
    // reg [31:0] Inst_Mem [INST_NUM - 1:0];

    
    always @(PC_Reg) begin
        Instruction = 0;
        case (PC_Reg[31:2])
            0: Instruction = 32'b1110_00_1_1101_0_0000_0000_000000010100; //MOV R0 ,#20 //R0 = 20
            1: Instruction = 32'b1110_00_1_1101_0_0000_0001_101000000001; //MOV R1 ,#4096 //R1 = 4096
            2: Instruction = 32'b1110_00_1_1101_0_0000_0010_000100000011; //MOV R2 ,#0xC0000000 //R2 = -1073741824
            3: Instruction = 32'b1110_00_0_0100_1_0010_0011_000000000010; //ADDS R3 ,R2,R2 //R3 = -2147483648 
            4: Instruction = 32'b1110_00_0_0101_0_0000_0100_000000000000; //ADC R4 ,R0,R0 //R4 = 41
            5: Instruction = 32'b1110_00_0_0010_0_0100_0101_000100000100; //SUB R5 ,R4,R4,LSL #2 //R5 = -123
            6: Instruction = 32'b1110_00_0_0110_0_0000_0110_000010100000; //SBC R6 ,R0,R0,LSR #1 //R6 = 10
            7: Instruction = 32'b1110_00_0_1100_0_0101_0111_000101000010; //ORR R7 ,R5,R2,ASR #2 //R7 = -123
            8: Instruction = 32'b1110_00_0_0000_0_0111_1000_000000000011; //AND R8 ,R7,R3 //R8 = -2147483648
            9: Instruction = 32'b1110_00_0_1111_0_0000_1001_000000000110; //MVN R9 ,R6 //R9 = -11
            10: Instruction = 32'b1110_00_0_0001_0_0100_1010_000000000101; //EOR R10,R4,R5 //R10 = -84
            11: Instruction = 32'b1110_00_0_1010_1_1000_0000_000000000110; //CMP R8 ,R6
            12: Instruction = 32'b0001_00_0_0100_0_0001_0001_000000000001; //ADDNE R1 ,R1,R1 //R1 = 8192
            13: Instruction = 32'b1110_00_0_1000_1_1001_0000_000000001000; //TST R9 ,R8
            14: Instruction = 32'b0000_00_0_0100_0_0010_0010_000000000010; //ADDEQ R2 ,R2,R2 //R2 = -1073741824
            15: Instruction = 32'b1110_00_1_1101_0_0000_0000_101100000001; //MOV R0 ,#1024
            16: Instruction = 32'b1110_01_0_0100_0_0000_0001_000000000000; //STR R1 ,[R0],#0 //MEM[1024] = 8192
            17: Instruction = 32'b1110_01_0_0100_1_0000_1011_000000000000; //LDR R11,[R0],#0 //R11 = 8192
            18: Instruction = 32'b1110_01_0_0100_0_0000_0010_000000000100; //STR R2 ,[R0],#4 //MEM[1028] = -1073741824
            19: Instruction = 32'b1110_01_0_0100_0_0000_0011_000000001000; //STR R3 ,[R0],#8 //MEM[1032] = -2147483648
            20: Instruction = 32'b1110_01_0_0100_0_0000_0100_000000001101; //STR R4 ,[R0],#13 //MEM[1036] = 41
            21: Instruction = 32'b1110_01_0_0100_0_0000_0101_000000010000; //STR R5 ,[R0],#16 //MEM[1040] = -123
            22: Instruction = 32'b1110_01_0_0100_0_0000_0110_000000010100; //STR R6 ,[R0],#20 //MEM[1044] = 10
            23: Instruction = 32'b1110_01_0_0100_1_0000_1010_000000000100; //LDR R10,[R0],#4 //R10 = -1073741824
            24: Instruction = 32'b1110_01_0_0100_0_0000_0111_000000011000; //STR R7 ,[R0],#24 //MEM[1048] = -123
            25: Instruction = 32'b1110_00_1_1101_0_0000_0001_000000000100; //MOV R1 ,#4 //R1 = 4
            26: Instruction = 32'b1110_00_1_1101_0_0000_0010_000000000000; //MOV R2 ,#0 //R2 = 0
            27: Instruction = 32'b1110_00_1_1101_0_0000_0011_000000000000; //MOV R3 ,#0 //R3 = 0
            28: Instruction = 32'b1110_00_0_0100_0_0000_0100_000100000011; //ADD R4 ,R0,R3,LSL #2
            29: Instruction = 32'b1110_01_0_0100_1_0100_0101_000000000000; //LDR R5 ,[R4],#0
            30: Instruction = 32'b1110_01_0_0100_1_0100_0110_000000000100; //LDR R6 ,[R4],#4
            31: Instruction = 32'b1110_00_0_1010_1_0101_0000_000000000110; //CMP R5 ,R6
            32: Instruction = 32'b1100_01_0_0100_0_0100_0110_000000000000; //STRGT R6 ,[R4],#0
            33: Instruction = 32'b1100_01_0_0100_0_0100_0101_000000000100; //STRGT R5 ,[R4],#4
            34: Instruction = 32'b1110_00_1_0100_0_0011_0011_000000000001; //ADD R3 ,R3,#1
            35: Instruction = 32'b1110_00_1_1010_1_0011_0000_000000000011; //CMP R3 ,#3
            36: Instruction = 32'b1011_10_1_0_111111111111111111110111 ; //BLT #-9
            37: Instruction = 32'b1110_00_1_0100_0_0010_0010_000000000001; //ADD R2 ,R2,#1
            38: Instruction = 32'b1110_00_0_1010_1_0010_0000_000000000001; //CMP R2 ,R1
            39: Instruction = 32'b1011_10_1_0_111111111111111111110011 ; //BLT #-13
            40: Instruction = 32'b1110_01_0_0100_1_0000_0001_000000000000; //LDR R1 ,[R0],#0 //R1 = -2147483648
            41: Instruction = 32'b1110_01_0_0100_1_0000_0010_000000000100; //LDR R2 ,[R0],#4 //R2 = -1073741824
            42: Instruction = 32'b1110_01_0_0100_1_0000_0011_000000001000; //LDR R3 ,[R0],#8 //R3 = 41
            43: Instruction = 32'b1110_01_0_0100_1_0000_0100_000000001100; //LDR R4 ,[R0],#12 //R4 = 8192
            44: Instruction = 32'b1110_01_0_0100_1_0000_0101_000000010000; //LDR R5 ,[R0],#16 //R5 = -123
            45: Instruction = 32'b1110_01_0_0100_1_0000_0110_000000010100; //LDR R6 ,[R0],#20 //R4 = 10
            46: Instruction = 32'b1110_10_1_0_111111111111111111111111 ; //B #-1

            default Instruction = {4'b1110, 28'b0};
        endcase
        
    end

    //PC_Reg
    always @(posedge clk, posedge rst) begin
        if(rst)
            PC_Reg <= 0;
        else if(~freeze)
            PC_Reg <= PC_In;
    end

    assign PC_In = Branch_taken ? BranchAddr : PC;
    assign PC = PC_Reg + 4;
    // assign Instruction = Inst_Mem[PC_Reg[$clog2(INST_NUM)+2:2]];
    
    

    
endmodule